module TwosToSignMag;

endmodule

module FloatingPointConvert;

endmodule

module Rounding;

endmodule